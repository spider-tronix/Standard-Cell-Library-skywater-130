.option scale=1E-6
.include "O:/sky130_fd_pr/models/r+c/res_typical__cap_typical__lin.spice"
.include "O:/sky130_fd_pr/models/r+c/res_typical__cap_typical.spice"
.include "O:/sky130_fd_pr/models/corners/tt.spice"

X1 Vdd A1 P001 N001 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X2 P001 A2 P002 N003 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X3 P002 A3 Y N004 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X4 Vdd B1 Y N002 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X5 Y B1 N006 N005 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X7 N006 A1 0 N007 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X8 N006 A2 0 N008 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X9 N006 A3 0 N009 sky130_fd_pr__nfet_01v8 l=0.18 w=2

V1 A1 0 PULSE(0 1.8 0 0 0 5 10)
V2 A2 0 0
V3 A3 0 0
V4 Vdd 0 1.8
V6 B1 0 1.8

.tran 0.001 50
.end