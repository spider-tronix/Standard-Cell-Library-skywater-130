.inc /home/akil/Skywater130spice/sky130.lib
M1 N004 A N007 N005 cmosn l=0.13u w=0.13u
M2 Vdd A N004 N002 cmosp l=0.13u w=0.13u
V1 Vdd 0 1.8
V2 A 0 PULSE(0 1.8 0 0 0 5 10)
M3 N007 B 0 N008 cmosn l=0.13u w=0.13u
M4 Vdd B N004 N003 cmosp l=0.13u w=0.13u
V3 B 0 1.8
M5 Y N004 0 N006 cmosn l=0.13u w=0.13u
M6 Vdd N004 Y N001 cmosp l=0.13u w=0.13u
.tran 10u 50
.end
