.option scale=1E-6
.include "O:/sky130_fd_pr/models/r+c/res_typical__cap_typical__lin.spice"
.include "O:/sky130_fd_pr/models/r+c/res_typical__cap_typical.spice"
.include "O:/sky130_fd_pr/models/corners/tt.spice"
X1 Vdd A1 P001 NC_01 sky130_fd_pr__pfet_01v8 l=0.18 w=1
X2 P001 A2 P002 N001 sky130_fd_pr__pfet_01v8 l=0.18 w=1
X3 P002 A3 P003 N003 sky130_fd_pr__pfet_01v8 l=0.18 w=1
X4 P003 A4 Y N004 sky130_fd_pr__pfet_01v8 l=0.18 w=1
X5 Vdd B1 Y N002 sky130_fd_pr__pfet_01v8 l=0.18 w=1
X6 Y B1 N006 N005 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X7 N006 A1 0 N007 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X8 N006 A2 0 N008 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X9 N006 A3 0 N009 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X10 N006 A4 0 N010 sky130_fd_pr__nfet_01v8 l=0.18 w=1
.end
