.option scale=1E-6
.include "/home/akil/sky130_fd_pr/models/r+c/res_typical__cap_typical__lin.spice"
.include "/home/akil/sky130_fd_pr/models/r+c/res_typical__cap_typical.spice"
.include "/home/akil/sky130_fd_pr/models/corners/tt.spice"

X1 Vdd N007 Y Vdd sky130_fd_pr__pfet_01v8 l=0.18 w=2
X2 Y N007 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X3 Vdd A N001 Vdd sky130_fd_pr__pfet_01v8 l=0.18 w=2
X4 Vdd B N001 Vdd sky130_fd_pr__pfet_01v8 l=0.18 w=2
X5 N001 A N002 N001 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X6 N001 C N002 N001 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X7 N002 B N007 N002 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X8 N002 C N007 N002 sky130_fd_pr__pfet_01v8 l=0.18 w=2
X9 N007 A N003 N003 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X10 N007 A N004 N004 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X11 N007 B N005 N005 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X12 N003 B 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X13 N004 C 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=2
X14 N005 C 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=2

CL Y 0 0.6pF
V1 A 0 PULSE(0 1.8 0 0.06n 0.06n 10.0n 20n)
V2 B 0 0
V3 C 0 1.8
V4 Vdd 0 1.8
.tran 0.1n 100n 
.end