* O:\VSD Intern\LT spice\Schematics\NAND.asc
M1 Y A N004 N003 cmosn l=0.13u w=2u
M2 Vdd A Y N001 cmosp l=0.13u w=2u
V1 Vdd 0 1.8
V2 A 0 PULSE(0 1.8 0 0 0 5n 10n)
M3 N004 B 0 N005 cmosn l=0.13u w=2u
M4 Vdd B Y N002 cmosp l=0.13u w=2u
V3 B 0 1.8
.tran 0.01n 50n
.model cmosn NMOS(
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.255e-06 wmax = 1.265e-06
+ level = 54
+ tnom = 30
+ version = 4.5
+ toxm = 4.148e-009
+ xj = 1.5e-007
+ lln = 1
+ lwn = 1
+ wln = 1
+ wwn = 1
+ lint = 1.1932e-008+0.0
+ ll = 0
+ lw = 0
+ lwl = 0
+ wint = 2.1859e-008+0.0
+ wl = 0
+ ww = 0
+ wwl = 0
+ xl = 0
+ xw = 0
+ mobmod = 0
+ binunit = 2
+ dwg = 0
+ dwb = 0
+ igcmod = 0
+ igbmod = 0
+ rgatemod = 0
+ rbodymod = 1
+ trnqsmod = 0
+ acnqsmod = 0
+ fnoimod = 1
+ tnoimod = 1
+ permod = 1
+ geomod = 0
+ rdsmod = 0
+ tempmod = 0
+ lintnoi = -1.0e-07
+ vfbsdoff = 0
+ lambda = 0
+ vtl = 0
+ lc = 5e-009
+ xn = 3
+ rnoia = 0.94
+ rnoib = 0.26
+ tnoia = 1.5e7
+ tnoib = 9.9e6
+ epsrox = 3.9
+ toxe = 4.148e-009
+ dtox = 0
+ ndep = 1.7e+017
+ nsd = 1e+020
+ rshg = 0.1
+ rsh = 1
+ vth0 = 0.49439+0.0
+ k1 = 0.90707349
+ k2 = -0.12949+0.0
+ k3 = 2
+ dvt0 = 0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600
+ dvt2w = 0.068
+ w0 = 0
+ k3b = 0.54
+ phin = 0
+ lpe0 = 1.0325e-007
+ lpeb = -7.082e-008
+ vbm = -3
+ dvtp0 = 0
+ dvtp1 = 0
+ vsat = 176320+0.0
+ ua = -1.1926e-009+0.0
+ ub = 2.1846e-018+0.0
+ uc = 8.1022e-011
+ rdsw = 65.968+0.0
+ prwb = 0
+ prwg = 0.021507
+ wr = 1
+ u0 = 0.030197+0.0
+ a0 = 1.5+0.0
+ keta = 0+0.0
+ a1 = 0
+ a2 = 0.42385546
+ ags = 1.25+0.0
+ b0 = 0+0.0
+ b1 = 0+0.0
+ eu = 1.67
+ rdswmin = 0
+ rdw = 0
+ rdwmin = 0
+ rsw = 0
+ rswmin = 0
+ voff = -0.20753+0.0
+ nfactor = 2.015+0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0+0.0
+ cit = 0
+ cdsc = 0
+ cdscb = 0
+ cdscd = 0.002052
+ eta0 = 0.00069413878+0.0
+ etab = -0.043998
+ dsub = 0.45862506
+ voffl = 5.8197729e-009
+ minv = 0
+ pclm = 0.14094+0.0
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 7.9141988e+008
+ pscbe2 = 1e-012
+ pvag = 0
+ delta = 0.01
+ alpha0 = 3e-008
+ alpha1 = 0.85
+ beta0 = 13.85
+ fprout = 0
+ pdits = 0+0.0
+ pditsl = 0
+ pditsd = 0+0.0
+ agidl = 0
+ bgidl = 2.3e+009
+ cgidl = 0.5
+ egidl = 0.8
+ aigbacc = 1
+ bigbacc = 0
+ cigbacc = 0
+ nigbacc = 0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0
+ poxedge = 1
+ pigcd = 1
+ ntox = 1
+ toxref = 4.148e-009
+ kt1 = -0.22096074+0.0
+ kt2 = -0.028878939
+ at = 40720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-011
+ ub1 = 7.0775317e-019
+ uc1 = 1.4718625e-010
+ kt1l = 0
+ prt = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbdb = 50
+ rbsb = 50
+ gbmin = 1e-012
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000E+07
+ af = 1
+ ef = 0.84
+ kf = 0
+ ntnoi = 1
+ dmcg = 0
+ dmcgt = 0
+ dmdg = 0
+ xgw = 0
+ xgl = 0
+ ngcon = 1
+ diomod = 1
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6e-10
+ xtis = 2
+ bvs = 11.7
+ xjbvs = 1
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
+ tpb = 0.0012287
+ tpbsw = 0
+ tpbswg = 0
+ tcj = 0.000792
+ tcjsw = 1e-005
+ tcjswg = 0
+ cgdo = 2.54e-010
+ cgso = 2.54e-010
+ cgbo = 1e-013
+ capmod = 2
+ xpart = 0
+ cgsl = 0
+ cgdl = 0
+ cf = 1.4067e-012
+ clc = 1e-007
+ cle = 0.6
+ dlc = 1.0494e-008+0.0+0.0
+ dwc = 0+0.0
+ vfbcv = -1
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
+ ngate = 1e+023
+ lwc = 0
+ llc = 0
+ lwlc = 0
+ wlc = 0
+ wwc = 0
+ wwlc = 0
+ ckappas = 0.6
+ cjs = 0.0013459
+ mjs = 0.44
+ pbs = 0.729
+ cjsws = 3.6001e-011
+ mjsws = 0.0009
+ pbsws = 0.2
+ cjswgs = 2.3347e-010
+ mjswgs = 0.8000
+ pbswgs = 0.95578
+ saref = 1.04e-06
+ sbref = 1.04e-06
+ wlod = 0
+ kvth0 = 9.8e-9
+ lkvth0 = 0
+ wkvth0 = 0.2e-6
+ pkvth0 = 0
+ llodvth = 0
+ wlodvth = 1
+ stk2 = 0
+ lodk2 = 1
+ lodeta0 = 1
+ ku0 = -2.7e-08
+ lku0 = 0
+ wku0 = 0
+ pku0 = 0
+ llodku0 = 0
+ wlodku0 = 1
+ kvsat = 0.2
+ steta0 = 0
+ tku0 = 0
+)
.model cmosp PMOS (
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.255e-06 wmax = 1.265e-06
+ level = 54
+ tnom = 30
+ version = 4.5
+ toxm = 4.23e-009
+ xj = 1.5e-007
+ lln = 1
+ lwn = 1
+ wln = 1
+ wwn = 1
+ lint = -1.3994e-008+0.0
+ ll = 0
+ lw = 0
+ lwl = 0
+ wint = 7.3039e-009+0.0
+ wl = 0
+ ww = 0
+ wwl = 0
+ xl = 0
+ xw = 0
+ mobmod = 0
+ binunit = 2
+ dwg = -5.722e-009
+ dwb = -1.7864e-008
+ igcmod = 0
+ igbmod = 0
+ rgatemod = 0
+ rbodymod = 1
+ trnqsmod = 0
+ acnqsmod = 0
+ fnoimod = 1
+ tnoimod = 1
+ permod = 1
+ geomod = 0
+ rdsmod = 0
+ tempmod = 0
+ lintnoi = -2.0e-07
+ vfbsdoff = 0
+ lambda = 0
+ vtl = 0
+ lc = 5e-009
+ xn = 3
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25e6
+ tnoib = 0.0e-6
+ epsrox = 3.9
+ toxe = 4.23e-009
+ dtox = 0
+ ndep = 1.7e+017
+ nsd = 1e+020
+ rshg = 0.1
+ rsh = 1
+ vth0 = -1.0652+0.0
+ k1 = 1.3152469
+ k2 = -0.27798063+0.0
+ k3 = -15.845
+ dvt0 = 4.4955
+ dvt1 = 0.294
+ dvt2 = 0.015
+ dvt0w = -4.9772
+ dvt1w = 1147200
+ dvt2w = -0.00896
+ w0 = 0
+ k3b = 2
+ phin = 0
+ lpe0 = 0
+ lpeb = 0
+ vbm = -3
+ dvtp0 = 0
+ dvtp1 = 0
+ vsat = 68611+0.0
+ ua = -2.4423e-009+0.0
+ ub = 2.0699352e-018+0.0
+ uc = 1.6133739e-013
+ rdsw = 547.88+0.0
+ prwb = -0.32348
+ prwg = 0.1376
+ wr = 1
+ u0 = 0.0025134+0.0
+ a0 = 0.91285081+0.0
+ keta = -0.020464881+0.0
+ a1 = 0
+ a2 = 0.87366558
+ ags = 1.25+0.0
+ b0 = 0+0.0
+ b1 = 0+0.0
+ eu = 1.67
+ rdswmin = 0
+ rdw = 0
+ rdwmin = 0
+ rsw = 0
+ rswmin = 0
+ voff = -0.25076476+0.0
+ nfactor = 1.9+0.0
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0+0.0
+ cit = 1e-005
+ cdsc = 0.00013
+ cdscb = 0.00078
+ cdscd = 0
+ eta0 = 0.21064695+0.0
+ etab = -0.014728557
+ dsub = 0.26
+ voffl = 0
+ minv = 0
+ pclm = 0.61630162+0.0
+ pdiblc1 = 0.14215108
+ pdiblc2 = 0.0026509038
+ pdiblcb = -0.15188768
+ drout = 1
+ pscbe1 = 8e+008
+ pscbe2 = 9.1788025e-009
+ pvag = 0
+ delta = 0.01
+ alpha0 = 1e-010
+ alpha1 = 1e-010
+ beta0 = 7.9381315
+ fprout = 0
+ pdits = 0+0.0
+ pditsl = 0
+ pditsd = 0+0.0
+ agidl = 4.0078966e-010+0.0
+ bgidl = 1e009+0.0
+ cgidl = 300+0.0
+ egidl = 0.1
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0
+ poxedge = 1
+ pigcd = 1
+ ntox = 1
+ toxref = 4.23e-009
+ kt1 = -0.70976+0.0
+ kt2 = -0.12
+ at = 50942
+ ute = -0.21243
+ ua1 = 1.8303e-010
+ ub1 = 3.6891e-019
+ uc1 = 6.4484e-012
+ kt1l = 0
+ prt = 0
+ xrcrg1 = 12
+ xrcrg2 = 1
+ rbpb = 50
+ rbpd = 50
+ rbps = 50
+ rbdb = 50
+ rbsb = 50
+ gbmin = 1e-012
+ noia = 1.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000E+07
+ af = 1
+ ef = 1.0
+ kf = 0
+ ntnoi = 1
+ dmcg = 0
+ dmcgt = 0
+ dmdg = 0
+ xgw = 0
+ xgl = 0
+ ngcon = 1
+ diomod = 1
+ njs = 1.3632
+ jss = 2.1483e-05
+ jsws = 8.040000000000001e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
+ tpb = 0.0020386
+ tpbsw = 0.001246
+ tpbswg = 0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2e-012
+ cgdo = 5.5e-11
+ cgso = 5.5e-11
+ cgbo = 0
+ capmod = 2
+ xpart = 0
+ cgsl = 1.0005e-011
+ cgdl = 1.0005e-011
+ cf = 1.2e-011
+ clc = 1e-007
+ cle = 0.6
+ dlc = -3e-09+0.0+0.0
+ dwc = 0+0.0
+ vfbcv = -0.14469
+ acde = 0.8
+ moin = 18.13
+ noff = 3.9
+ voffcv = -0.10701
+ ngate = 1e+023
+ lwc = 0
+ llc = 0
+ lwlc = 0
+ wlc = 0
+ wwc = 0
+ wwlc = 0
+ ckappas = 0.6
+ cjs = 0.00074079
+ mjs = 0.34629
+ pbs = 0.6587
+ cjsws = 9.88e-011
+ mjsws = 0.29781
+ pbsws = 0.7418
+ cjswgs = 2.3894e-010
+ mjswgs = 0.9274
+ pbswgs = 1.4338
+ saref = 1.04e-06
+ sbref = 1.04e-06
+ wlod = 0+0.0
+ kvth0 = 0+0.0
+ lkvth0 = 0+0.0
+ wkvth0 = 0+0.0
+ pkvth0 = 0
+ llodvth = 0
+ wlodvth = 1
+ stk2 = 0
+ lodk2 = 1
+ lodeta0 = 1
+ ku0 = 0+0.0
+ lku0 = 0+0.0
+ wku0 = 0+0.0
+ pku0 = 0
+ llodku0 = 0
+ wlodku0 = 1
+ kvsat = 0+0.0
+ steta0 = 0
+ tku0 = 0
+)
.end
