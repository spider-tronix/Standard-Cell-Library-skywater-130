.option scale=1E-6
.include "/home/akil/sky130_fd_pr/models/r+c/res_typical__cap_typical__lin.spice"
.include "/home/akil/sky130_fd_pr/models/r+c/res_typical__cap_typical.spice"
.include "/home/akil/sky130_fd_pr/models/corners/tt.spice"

X1 Vdd A1 N001 Vdd sky130_fd_pr__pfet_01v8 l=0.18 w=4.6
X2 N001 A2 N002 N001 sky130_fd_pr__pfet_01v8 l=0.18 w=4.6
X3 N002 A3 N003 N002 sky130_fd_pr__pfet_01v8 l=0.18 w=4.6
X4 N003 A4 Y N003 sky130_fd_pr__pfet_01v8 l=0.18 w=4.6
X5 Vdd B1 Y Vdd sky130_fd_pr__pfet_01v8 l=0.18 w=1
X6 Y B1 N004 N004 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X7 N004 A1 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X8 N004 A2 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X9 N004 A3 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=1
X10 N004 A4 0 0 sky130_fd_pr__nfet_01v8 l=0.18 w=1

CL Y 0 0.6pF

V1 A1 0 PULSE(0 1.8 0 0.06n 0.06n 10.0n 20n)
V2 A2 0 0
V3 A3 0 0
V4 Vdd 0 1.8
V5 B1 0 1.8
V6 A4 0 0

.tran 0.1n 100n
.end